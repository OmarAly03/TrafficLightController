library verilog;
use verilog.vl_types.all;
entity TLC_Project_vlg_vec_tst is
end TLC_Project_vlg_vec_tst;
